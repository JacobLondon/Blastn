library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

entity Top is
    port (
        clk : in  STD_LOGIC;
        rst : in  STD_LOGIC;
        rx  : in  STD_LOGIC;
        tx  : out STD_LOGIC
    );
end Top;

architecture Blastn of Top is
    
    
    
begin

    

end Blastn;
